From Stdlib Require Import Utf8 ZArith.
From Crypto Require Import Sigma  Elgamal.
From Utility Require Import Zpstar Util.
From Frontend Require Import Approval.
From Backend Require Import HeliosTally.
From Examples Require Import primeP primeQ. 
Import Vspace Schnorr Zpfield Zpgroup.

(* 2024 https://vote.heliosvoting.org/helios/elections/a447fe8a-80c8-11ef-923c-7aae6cdba09d *)
(* 2023 https://vote.heliosvoting.org/helios/elections/c3dd2456-6a89-11ee-b981-bad8622d1122 *)
(* 2022 https://vote.heliosvoting.org/helios/elections/2565efe0-4958-11ed-b89e-7ad723fa8d9f *)
(* 
    In all these elections, p, q, and g are the same but h is different.
    We create a module Helios to encapsulate these parameters and the function to compute final count.
    In Helios, we create a sub-module IACR2022, IACR2023, IACR2024 for each year's election parameters
    and since only h is different, we define h separately in each sub-module.

*)
Section Helios.

  (* 256 bit Prime q*)
  Definition q : Z := 61329566248342901292543872769978950870633559608669337131139375508370458778917%Z.
  (* Eval compute in  N.size 61329566248342901292543872769978950870633559608669337131139375508370458778917. *)

  Theorem prime_q : Znumtheory.prime q.
  Proof.
  Admitted.

  (* 2048 bit Prime p *)
  Definition p : Z := 16328632084933010002384055033805457329601614771185955389739167309086214800406465799038583634953752941675645562182498120750264980492381375579367675648771293800310370964745767014243638518442553823973482995267304044326777047662957480269391322789378384619428596446446984694306187644767462460965622580087564339212631775817895958409016676398975671266179637898557687317076177218843233150695157881061257053019133078545928983562221396313169622475509818442661047018436264806901023966236718367204710755935899013750306107738002364137917426595737403871114187750804346564731250609196846638183903982387884578266136503697493474682071%Z.

  Theorem prime_p : Znumtheory.prime p.
  Proof.
  Admitted.
  
  (* 
  Eval compute in N.size 16328632084933010002384055033805457329601614771185955389739167309086214800406465799038583634953752941675645562182498120750264980492381375579367675648771293800310370964745767014243638518442553823973482995267304044326777047662957480269391322789378384619428596446446984694306187644767462460965622580087564339212631775817895958409016676398975671266179637898557687317076177218843233150695157881061257053019133078545928983562221396313169622475509818442661047018436264806901023966236718367204710755935899013750306107738002364137917426595737403871114187750804346564731250609196846638183903982387884578266136503697493474682071.
  *)
  

  
  (* safe prime *)
  Definition k : Z := Z.div p q. 

  Theorem safe_prime : p = (k * q + 1)%Z.
  Proof. vm_cast_no_check (eq_refl p).  Qed.

  Definition gval : Z := 14887492224963187634282421537186040801304008017743492304481737382571933937568724473847106029915040150784031882206090286938661464458896494215273989547889201144857352611058572236578734319505128042602372864570426550855201448111746579871811249114781674309062693442442368697449970648232621880001709535143047913661432883287150003429802392229361583608686643243349727791976247247948618930423866180410558458272606627111270040091203073580238905303994472202930783207472394578498507764703191288249547659899997131166130259700604433891232298182348403175947450284433411265966789131024573629546048637848902243503970966798589660808533%Z.

  
  Definition g : @Schnorr_group p q.
  Proof. 
    refine 
      {| Schnorr.v := gval;
      Ha := conj eq_refl eq_refl : (0 < gval < p)%Z;
      Hb := _ (* eq_refl : (Zpow_mod gval q p)%Z = 1%Z *)|}.
    vm_cast_no_check (eq_refl (Zpow_facts.Zpow_mod gval q p)). 
  Defined.

  (* 
  (* public key that changes each year *)
  Definition hval2024 : Z := 7046735122051745594868985795786176392951854019485729367165971776021501311096201521482383017242860186177215354508901537446984239682993203747271798136868016921883953390308299741287014686008274215001426444189972901892121945650333202105534018888882197552388434304153312708859768386971193915314738375008791798536164901595463713712574129466783480981077498017586306273866594394401039338841105927980179401433149438028686338492134818995843560711439253445043076178166622915392760675509176356257990398772342230639242314592068285808565623831103115873314006496120730338309413064358649726464219249576117734308027594482849210379533%Z. 

  (* 2024 election had 7 candidates. *)
  Definition h2024 : @Schnorr_group p q. 
  Proof. 
    refine
    {| 
      Schnorr.v := hval2024;
      Ha := conj eq_refl eq_refl : (0 < hval2024 < p)%Z;
      Hb := _ (* eq_refl : (Zpow_mod gval q p)%Z = 1%Z *)|}.
      vm_cast_no_check (eq_refl (Zpow_facts.Zpow_mod hval2024 q p)). 
  Defined.
  *)
  
  Definition hval2023 : Z := 
  13396065692002658190209213918774474470352093532579311681373807462187387355392940152980335043314279566135304465932321505117199458458691703887061297402530469179036279081346297942647302277396696748068899327427173907449796015294748375392495725034007822567958711624538227213705702406059840254658956003363562396354441345335395156606116320333570202517406626946073836664803134614881201398731965680643717511846389946291487290758319833954626923013580650083154183407956145565561747950100196644243904999390949701945284494916708366378558442200750198240994823297922478004889699261017557130340798590600460133638817687107827197373627%Z. 

  (* 2023 election had 6 candidates. *)
  Definition h2023 : @Schnorr_group p q.
  Proof. 
    refine
    {| 
      Schnorr.v := hval2023;
      Ha := conj eq_refl eq_refl : (0 < hval2023 < p)%Z;
      Hb := _ (* eq_refl : (Zpow_mod gval q p)%Z = 1%Z *)|}.
      vm_cast_no_check (eq_refl (Zpow_facts.Zpow_mod hval2023 q p)). 
  Defined.

  (*
  Definition hval2022 : Z := 8104845379024737751179395306670759432773921014970882975863017259159755939139951543095628383118775025713998854402843031464380570059038830419901388411272123087558933778250276505787888006021311325046668471999761357537697020047483370216202604781057219914810417006866960196819046287455995543070553744002406912570654087687482296200647340672422169310090868180700021366750036313854837787159248832939897674578629261242593839595526247341093517097574130759323514013160719386447363900873086825944386111943104164303052321342357566387615463613007214084782471120717452853735668684321143425769815893710067621236208575779675723538479%Z.

  (* 2022 election had 6 candidates. *)
  Definition h2022 : @Schnorr_group p q.
  Proof. 
    refine
    {| 
      Schnorr.v := hval2022;
      Ha := conj eq_refl eq_refl : (0 < hval2022 < p)%Z;
      Hb := _ (* eq_refl : (Zpow_mod gval q p)%Z = 1%Z *)|}.
      vm_cast_no_check (eq_refl (Zpow_facts.Zpow_mod hval2022 q p)). 
  Defined.

  *)

  (* enc of public key that changes each year *)

  

  Definition compute_final_count_ins {n m : nat} (h : @Schnorr_group p q)
    (bs : list (@ballot (@Zp q) (@Schnorr_group p q) n)) 
    (ts : Vector.t (@tallier (@Zp q) (@Schnorr_group p q) n) (1 + m))
    (pt : Vector.t (@Zp q) n) : 
    existsT (bfinal : bool) 
    (vbs inbs : list (@ballot (@Zp q) (@Schnorr_group p q) n)),
    @count (@Zp q)  
    (@Zpfield.zero q prime_q) 
    (@Zpfield.one q prime_q) zp_add zp_dec 
    (@Schnorr_group p q)  (@Schnorr.one p q prime_p prime_q)
    (@inv_schnorr_group _ p q safe_prime prime_p prime_q)
    (@mul_schnorr_group p q prime_p prime_q)
    (@pow k p q safe_prime prime_p prime_q)
    Schnorr.dec_zpstar n m g h  
    (finished bs vbs inbs ts pt bfinal).
  Proof.
    refine(@compute_final_count (@Zp q) 
    (@Zpfield.zero q prime_q) 
    (@Zpfield.one q prime_q) zp_add zp_dec 
    (@Schnorr_group p q) (@Schnorr.one p q prime_p prime_q)
    (@inv_schnorr_group _ p q safe_prime prime_p prime_q)
    (@mul_schnorr_group p q prime_p prime_q)
    (@pow k p q safe_prime prime_p prime_q)
    Schnorr.dec_zpstar n m g h bs ts pt).
  Defined.

End Helios.

  